module nand_gate(
  input a,b,
  output out);

  nand(out,a,b);

endmodule
