module nor_gate(
  input a, b,
  output out);

  nor(out,a,b);

endmodule
