module simple_alu(
  input [3:0]a,b,
  input [2:0]sel,
  output reg [3:0]result,
  output reg carry);

  always @(*) begin
  case(sel)
   3'b000 : {carry,result} = a+b;
   3'b001 : {carry,result} = a-b;
   3'b010 : result = a&b;
   3'b011 : result = a|b;
   3'b100 : result = a^b;
   3'b101 : result = a~^b;
   3'b110 : result = a/b;
   3'b111 : result = a%b;
   default : result = 4'b0000;
  endcase
  end
endmodule
