module dff_async_reset(
    input clk,
    input reset,
    input d,
    output reg q);
    always @(posedge clk or posedge reset) begin
        if (reset)
            q <= 1'b0;
        else
            q <= d;
end
endmodule
