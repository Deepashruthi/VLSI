module portdeclaration_pre2001(y,a,b);
   input a,b;
   output y;
   assign y=a&b;
endmodule
