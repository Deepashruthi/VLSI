module portdeclaration_post2001(output y,input a,b);
   assign y=a&b;
endmodule
